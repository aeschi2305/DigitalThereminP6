-- altera vhdl_input_version vhdl_2008
-----------------------------------------------------
-- Project : Digital Theremin
-----------------------------------------------------
-- File    : FIR_Decimation.vhd
-- Author  : dennis.aeschbacher@students.fhnw.ch
-----------------------------------------------------
-- Description : Applies an FIR Filter and Decimates the sampling Frequency by the factor dec
-----------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity fir_filter_pitch is
generic (
    N : natural := 13; --Number of Filter Coefficients
    M : natural := 29; --Number of Input Bits
    O : natural := 27 --Number of Output Bits
);
port (
  clk        : in  std_ulogic;
  reset_n       : in  std_ulogic;
  en_in        : in boolean;                  -- input enable
  en_out       : out std_ulogic;                 -- output enable
  en_out_dec   : out std_ulogic;                 -- output enable decimation
  i_data       : in  signed( M-1 downto 0);   -- data input
  o_data_dec   : out signed( O-1 downto 0);  -- data output
  o_data       : out signed( O-1 downto 0)  -- data output
);
end entity fir_filter_pitch;

architecture rtl of fir_filter_pitch is
type coeff_type is array (0 to N-1) of signed (O-1 downto 0);
constant addstages : natural := N-1; -- Number of summation stages
constant coeffs : coeff_type :=  ("000001101001110110111101",
                                  "000000101001101010011000",
                                  "000000110001001100111111",
                                  "000000111001000011011010",
                                  "000001000001001100101001",
                                  "000001001001100100000101",
                                  "000001010001111100001101",
                                  "000001011010010000010101",
                                  "000001100010010111100010",
                                  "000001101010001101110111",
                                  "000001110001100111110010",
                                  "000001111000011111011100",
                                  "000001111110101010001111",
                                  "000010000100000101001100",
                                  "000010001000101000011011",
                                  "000010001100010010010101",
                                  "000010001110111011101000",
                                  "000010010000100011110110",
                                  "000010010001000101110110",
                                  "000010010000100011110110",
                                  "000010001110111011101000",
                                  "000010001100010010010101",
                                  "000010001000101000011011",
                                  "000010000100000101001100",
                                  "000001111110101010001111",
                                  "000001111000011111011100",
                                  "000001110001100111110010",
                                  "000001101010001101110111",
                                  "000001100010010111100010",
                                  "000001011010010000010101",
                                  "000001010001111100001101",
                                  "000001001001100100000101",
                                  "000001000001001100101001",
                                  "000000111001000011011010",
                                  "000000110001001100111111",
                                  "000000101001101010011000",
                                  "000001101001110110111101");

type t_data_pipe      is array (0 to N-1) of signed(O-1  downto 0);
type t_mult           is array (0 to N-1) of signed(O*2-1    downto 0);
signal p_data_in_reg               : t_data_pipe;
signal p_data_in_cmb               : t_data_pipe;
signal p_data_out_reg              : signed(O-1 downto 0);
signal p_data_out_cmb              : signed(O-1 downto 0);

signal p_data_out_dec_reg              : signed(O-1 downto 0);

signal count_reg         : natural range 0 to 25;
signal count_cmb         : natural range 0 to 26;

begin

 p_reg : process(reset_n,clk)
    begin
        if reset_n = '0' then
            l_mult : for ii in 0 to N-1 loop
              p_data_in_reg(ii) <= (others => '0');
            end loop l_mult;
            p_data_out_reg <= (others => '0');
            en_out <= '0';
        elsif rising_edge(clk) then
            en_out <= '0';
            if en_in = true then 
              p_data_in_reg <= p_data_in_cmb;
              p_data_out_reg <= p_data_out_cmb;
              en_out <= '1';
            end if;
        end if;
    end process p_reg;

  p_reg_dec : process(reset_n,clk)
    begin
        if reset_n = '0' then
            
        elsif rising_edge(clk) then
            if count_reg = 24 then
              p_data_out_dec_reg <= p_data_out_reg;
              count_reg <= 0;
            else
              count_reg <= count_cmb;
            end if;
        end if;
    end process p_reg_dec;

p_cmb : process(all)
    variable mult   : t_mult;
    variable sum    : signed(O*2-1 downto 0);
      begin 
        p_data_in_cmb <= i_data(M-1 downto M-O) & p_data_in_reg(0 to p_data_in_reg'length-2);
        l_mult : for ii in 0 to N-1 loop
            mult(ii) := p_data_in_reg(ii)*coeffs(ii);
        end loop l_mult;
        sum := to_signed(0,sum'length);
        l_add : for ii in 0 to N-1 loop
            sum := sum+mult(ii);
        end loop l_add;
        p_data_out_cmb <= sum(O*2-1 downto O);
        
        count_cmb <= count_reg + 1;
    end process p_cmb;

    o_data <= p_data_out_reg; 
    o_data <= p_data_out_dec_reg; 
end rtl;