-- Test1kHz.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test1kHz is
	port (
		clk_clk                       : in    std_logic := '0'; --                   clk.clk
		codecdigitalinterface_BCLK    : in    std_logic := '0'; -- codecdigitalinterface.BCLK
		codecdigitalinterface_DACDAT  : out   std_logic;        --                      .DACDAT
		codecdigitalinterface_DACLRCK : in    std_logic := '0'; --                      .DACLRCK
		codeci2c_SDAT                 : inout std_logic := '0'; --              codeci2c.SDAT
		codeci2c_SCLK                 : out   std_logic;        --                      .SCLK
		reset_reset_n                 : in    std_logic := '0';  --                 reset.reset_n
		AUD_XCK           			  : out std_logic

	);
end entity Test1kHz;

architecture rtl of Test1kHz is
	component sine1kHz is
		generic (
			count_freq : integer := 47;
			count_samp : integer := 256
		);
		port (
			reset         : in  std_logic                     := 'X'; -- reset
			clk           : in  std_logic                     := 'X'; -- clk
			aso_seL_ready : in  std_logic                     := 'X'; -- ready
			aso_seL_valid : out std_logic;                            -- valid
			aso_seL_data  : out std_logic_vector(23 downto 0);        -- data
			aso_seR_ready : in  std_logic                     := 'X'; -- ready
			aso_seR_valid : out std_logic;                            -- valid
			aso_seR_data  : out std_logic_vector(23 downto 0)         -- data
		);
	end component sine1kHz;

	component Test1kHz_audio_0 is
		port (
			clk                          : in  std_logic                     := 'X';             -- clk
			reset                        : in  std_logic                     := 'X';             -- reset
	--		from_adc_left_channel_ready  : in  std_logic                     := 'X';             -- ready
	--		from_adc_left_channel_data   : out std_logic_vector(23 downto 0);                    -- data
	--		from_adc_left_channel_valid  : out std_logic;                                        -- valid
	--		from_adc_right_channel_ready : in  std_logic                     := 'X';             -- ready
	--		from_adc_right_channel_data  : out std_logic_vector(23 downto 0);                    -- data
	--		from_adc_right_channel_valid : out std_logic;                                        -- valid
			to_dac_left_channel_data     : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_left_channel_valid    : in  std_logic                     := 'X';             -- valid
			to_dac_left_channel_ready    : out std_logic;                                        -- ready
			to_dac_right_channel_data    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_dac_right_channel_valid   : in  std_logic                     := 'X';             -- valid
			to_dac_right_channel_ready   : out std_logic;                                        -- ready
			AUD_BCLK                     : in  std_logic                     := 'X';             -- export
			AUD_DACDAT                   : out std_logic;                                        -- export
			AUD_DACLRCK                  : in  std_logic                     := 'X'              -- export
		);
	end component Test1kHz_audio_0;

	component Test1kHz_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component Test1kHz_audio_and_video_config_0;

	component Test1kHz_audio_pll_0 is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			audio_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Test1kHz_audio_pll_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal test1khzsinecomponent_0_sel_valid : std_logic;                     -- Test1kHzSineComponent_0:aso_seL_valid -> audio_0:to_dac_left_channel_valid
	signal test1khzsinecomponent_0_sel_data  : std_logic_vector(23 downto 0); -- Test1kHzSineComponent_0:aso_seL_data -> audio_0:to_dac_left_channel_data
	signal test1khzsinecomponent_0_sel_ready : std_logic;                     -- audio_0:to_dac_left_channel_ready -> Test1kHzSineComponent_0:aso_seL_ready
	signal test1khzsinecomponent_0_ser_valid : std_logic;                     -- Test1kHzSineComponent_0:aso_seR_valid -> audio_0:to_dac_right_channel_valid
	signal test1khzsinecomponent_0_ser_data  : std_logic_vector(23 downto 0); -- Test1kHzSineComponent_0:aso_seR_data -> audio_0:to_dac_right_channel_data
	signal test1khzsinecomponent_0_ser_ready : std_logic;                     -- audio_0:to_dac_right_channel_ready -> Test1kHzSineComponent_0:aso_seR_ready
	signal audio_pll_0_audio_clk_clk         : std_logic;                     -- audio_pll_0:audio_clk_clk -> [Test1kHzSineComponent_0:clk, audio_0:clk, audio_and_video_config_0:clk, rst_controller:clk]
	signal rst_controller_reset_out_reset    : std_logic;                     -- rst_controller:reset_out -> [Test1kHzSineComponent_0:reset, audio_0:reset, audio_and_video_config_0:reset]
	signal audio_pll_0_reset_source_reset    : std_logic;                     -- audio_pll_0:reset_source_reset -> rst_controller:reset_in0
	signal reset_reset_n_ports_inv           : std_logic;                     -- reset_reset_n:inv -> audio_pll_0:ref_reset_reset

begin
	
	AUD_XCK <= audio_pll_0_audio_clk_clk;

	test1khzsinecomponent_0 : component sine1kHz
		generic map (
			count_freq => 47,
			count_samp => 256
		)
		port map (
			reset         => rst_controller_reset_out_reset,    -- reset.reset
			clk           => audio_pll_0_audio_clk_clk,         -- clock.clk
			aso_seL_ready => test1khzsinecomponent_0_sel_ready, --   sel.ready
			aso_seL_valid => test1khzsinecomponent_0_sel_valid, --      .valid
			aso_seL_data  => test1khzsinecomponent_0_sel_data,  --      .data
			aso_seR_ready => test1khzsinecomponent_0_ser_ready, --   ser.ready
			aso_seR_valid => test1khzsinecomponent_0_ser_valid, --      .valid
			aso_seR_data  => test1khzsinecomponent_0_ser_data   --      .data
		);

	audio_0 : component Test1kHz_audio_0
		port map (
			clk                          => audio_pll_0_audio_clk_clk,         --                         clk.clk
			reset                        => rst_controller_reset_out_reset,    --                       reset.reset
	--		from_adc_left_channel_ready  => open,                              --  avalon_left_channel_source.ready
	--		from_adc_left_channel_data   => open,                              --                            .data
	--		from_adc_left_channel_valid  => open,                              --                            .valid
	--		from_adc_right_channel_ready => open,                              -- avalon_right_channel_source.ready
	--		from_adc_right_channel_data  => open,                              --                            .data
	--		from_adc_right_channel_valid => open,                              --                            .valid
			to_dac_left_channel_data     => test1khzsinecomponent_0_sel_data,  --    avalon_left_channel_sink.data
			to_dac_left_channel_valid    => test1khzsinecomponent_0_sel_valid, --                            .valid
			to_dac_left_channel_ready    => test1khzsinecomponent_0_sel_ready, --                            .ready
			to_dac_right_channel_data    => test1khzsinecomponent_0_ser_data,  --   avalon_right_channel_sink.data
			to_dac_right_channel_valid   => test1khzsinecomponent_0_ser_valid, --                            .valid
			to_dac_right_channel_ready   => test1khzsinecomponent_0_ser_ready, --                            .ready
			AUD_BCLK                     => codecdigitalinterface_BCLK,        --          external_interface.export
			AUD_DACDAT                   => codecdigitalinterface_DACDAT,      --                            .export
			AUD_DACLRCK                  => codecdigitalinterface_DACLRCK      --                            .export
		);

	audio_and_video_config_0 : component Test1kHz_audio_and_video_config_0
		port map (
			clk         => audio_pll_0_audio_clk_clk,      --                    clk.clk
			reset       => rst_controller_reset_out_reset, --                  reset.reset
			address     => open,                           -- avalon_av_config_slave.address
			byteenable  => open,                           --                       .byteenable
			read        => open,                           --                       .read
			write       => open,                           --                       .write
			writedata   => open,                           --                       .writedata
			readdata    => open,                           --                       .readdata
			waitrequest => open,                           --                       .waitrequest
			I2C_SDAT    => codeci2c_SDAT,                  --     external_interface.export
			I2C_SCLK    => codeci2c_SCLK                   --                       .export
		);

	audio_pll_0 : component Test1kHz_audio_pll_0
		port map (
			ref_clk_clk        => clk_clk,                        --      ref_clk.clk
			ref_reset_reset    => reset_reset_n_ports_inv,        --    ref_reset.reset
			audio_clk_clk      => audio_pll_0_audio_clk_clk,      --    audio_clk.clk
			reset_source_reset => audio_pll_0_reset_source_reset  -- reset_source.reset
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => audio_pll_0_reset_source_reset, -- reset_in0.reset
			clk            => audio_pll_0_audio_clk_clk,      --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of Test1kHz
