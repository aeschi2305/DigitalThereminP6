-- system.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system is
	port (
		aud_xck_clk                                      : out   std_logic;                                        --                                     aud_xck.clk
		audio_and_video_config_0_external_interface_SDAT : inout std_logic                     := '0';             -- audio_and_video_config_0_external_interface.SDAT
		audio_and_video_config_0_external_interface_SCLK : out   std_logic;                                        --                                            .SCLK
		bclk_export                                      : in    std_logic                     := '0';             --                                        bclk.export
		clk_clk                                          : in    std_logic                     := '0';             --                                         clk.clk
		dacdat_export                                    : out   std_logic;                                        --                                      dacdat.export
		daclrck_export                                   : in    std_logic                     := '0';             --                                     daclrck.export
		dram_ctrl_wire_addr                              : out   std_logic_vector(12 downto 0);                    --                              dram_ctrl_wire.addr
		dram_ctrl_wire_ba                                : out   std_logic_vector(1 downto 0);                     --                                            .ba
		dram_ctrl_wire_cas_n                             : out   std_logic;                                        --                                            .cas_n
		dram_ctrl_wire_cke                               : out   std_logic;                                        --                                            .cke
		dram_ctrl_wire_cs_n                              : out   std_logic;                                        --                                            .cs_n
		dram_ctrl_wire_dq                                : inout std_logic_vector(15 downto 0) := (others => '0'); --                                            .dq
		dram_ctrl_wire_dqm                               : out   std_logic_vector(1 downto 0);                     --                                            .dqm
		dram_ctrl_wire_ras_n                             : out   std_logic;                                        --                                            .ras_n
		dram_ctrl_wire_we_n                              : out   std_logic;                                        --                                            .we_n
		lcd_controller_conduit_end_lt24_cs               : out   std_logic;                                        --                  lcd_controller_conduit_end.lt24_cs
		lcd_controller_conduit_end_lt24_data             : out   std_logic_vector(15 downto 0);                    --                                            .lt24_data
		lcd_controller_conduit_end_lt24_rd               : out   std_logic;                                        --                                            .lt24_rd
		lcd_controller_conduit_end_lt24_wr               : out   std_logic;                                        --                                            .lt24_wr
		lcd_controller_conduit_end_lt24_rs               : out   std_logic;                                        --                                            .lt24_rs
		lcd_reset_n_external_connection_export           : out   std_logic;                                        --             lcd_reset_n_external_connection.export
		led_delay_export                                 : out   std_logic;                                        --                                   led_delay.export
		led_gli_export                                   : out   std_logic;                                        --                                     led_gli.export
		led_vol_export                                   : out   std_logic;                                        --                                     led_vol.export
		reset_reset_n                                    : in    std_logic                     := '0';             --                                       reset.reset_n
		sdram_clk_clk                                    : out   std_logic;                                        --                                   sdram_clk.clk
		touch_panel_busy_external_connection_export      : in    std_logic                     := '0';             --        touch_panel_busy_external_connection.export
		touch_panel_pen_irq_n_external_connection_export : in    std_logic                     := '0';             --   touch_panel_pen_irq_n_external_connection.export
		touch_panel_spi_external_MISO                    : in    std_logic                     := '0';             --                    touch_panel_spi_external.MISO
		touch_panel_spi_external_MOSI                    : out   std_logic;                                        --                                            .MOSI
		touch_panel_spi_external_SCLK                    : out   std_logic;                                        --                                            .SCLK
		touch_panel_spi_external_SS_n                    : out   std_logic                                         --                                            .SS_n
	);
end entity system;

architecture rtl of system is
	component LT24_Controller is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			reset_n        : in  std_logic                     := 'X';             -- reset_n
			s_chipselect_n : in  std_logic                     := 'X';             -- chipselect_n
			s_write_n      : in  std_logic                     := 'X';             -- write_n
			s_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s_address      : in  std_logic                     := 'X';             -- address
			lt24_cs        : out std_logic;                                        -- lt24_cs
			lt24_data      : out std_logic_vector(15 downto 0);                    -- lt24_data
			lt24_rd        : out std_logic;                                        -- lt24_rd
			lt24_wr        : out std_logic;                                        -- lt24_wr
			lt24_rs        : out std_logic                                         -- lt24_rs
		);
	end component LT24_Controller;

	component system_LCD_Reset_N is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component system_LCD_Reset_N;

	component pitch_dummy is
		generic (
			dat_len_avl : natural                       := 31;
			data_freq   : std_logic_vector(31 downto 0) := "00000000000000001111101000000000";
			data_freq1  : std_logic_vector(31 downto 0) := "00000000000000000111110100000000"
		);
		port (
			avs_sP_address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avs_sP_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			avs_sP_write     : in  std_logic                     := 'X';             -- write
			avs_sP_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			coe_led_gli      : out std_logic;                                        -- export
			rsi_reset_n      : in  std_logic                     := 'X';             -- reset_n
			csi_clk          : in  std_logic                     := 'X';             -- clk
			coe_led_delay    : out std_logic                                         -- export
		);
	end component pitch_dummy;

	component volume_dummy is
		generic (
			dat_len_avl : natural                       := 31;
			data_freq   : std_logic_vector(31 downto 0) := "00000000000000001111101000000000";
			data_freq1  : std_logic_vector(31 downto 0) := "00000000000000000111110100000000"
		);
		port (
			avs_sP_address   : in  std_logic                     := 'X';             -- address
			avs_sP_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			avs_sP_write     : in  std_logic                     := 'X';             -- write
			avs_sP_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			coe_led_vol      : out std_logic;                                        -- export
			rsi_reset_n      : in  std_logic                     := 'X';             -- reset_n
			csi_clk          : in  std_logic                     := 'X'              -- clk
		);
	end component volume_dummy;

	component system_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component system_audio_and_video_config_0;

	component system_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component system_cpu;

	component system_dram_ctrl is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_dram_ctrl;

	component system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_jtag_uart;

	component system_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			outclk_3 : out std_logic;        -- clk
			outclk_4 : out std_logic;        -- clk
			outclk_5 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component system_pll;

	component system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component system_sysid;

	component system_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component system_timer;

	component sine1kHz is
		port (
			reset_n          : in  std_logic := 'X'; -- reset_n
			clk              : in  std_logic := 'X'; -- clk
			coe_AUD2_DACDAT  : out std_logic;        -- export
			coe_AUD1_BCLK    : in  std_logic := 'X'; -- export
			coe_AUD3_DACLRCK : in  std_logic := 'X'  -- export
		);
	end component sine1kHz;

	component system_touch_panel_busy is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component system_touch_panel_busy;

	component system_touch_panel_pen_irq_n is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component system_touch_panel_pen_irq_n;

	component system_touch_panel_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component system_touch_panel_spi;

	component system_mm_interconnect_0 is
		port (
			pll_outclk0_clk                                             : in  std_logic                     := 'X';             -- clk
			pll_outclk1_clk                                             : in  std_logic                     := 'X';             -- clk
			pll_outclk3_clk                                             : in  std_logic                     := 'X';             -- clk
			audio_and_video_config_0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			cpu_reset_reset_bridge_in_reset_reset                       : in  std_logic                     := 'X';             -- reset
			dram_ctrl_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			LCD_Controller_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                     : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                 : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                        : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                    : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                               : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                       : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                 : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                              : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                          : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                 : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                        : out std_logic;                                        -- readdatavalid
			audio_and_video_config_0_avalon_av_config_slave_address     : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_0_avalon_av_config_slave_write       : out std_logic;                                        -- write
			audio_and_video_config_0_avalon_av_config_slave_read        : out std_logic;                                        -- read
			audio_and_video_config_0_avalon_av_config_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_address                                 : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                   : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                    : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                             : out std_logic;                                        -- debugaccess
			dram_ctrl_s1_address                                        : out std_logic_vector(24 downto 0);                    -- address
			dram_ctrl_s1_write                                          : out std_logic;                                        -- write
			dram_ctrl_s1_read                                           : out std_logic;                                        -- read
			dram_ctrl_s1_readdata                                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			dram_ctrl_s1_writedata                                      : out std_logic_vector(15 downto 0);                    -- writedata
			dram_ctrl_s1_byteenable                                     : out std_logic_vector(1 downto 0);                     -- byteenable
			dram_ctrl_s1_readdatavalid                                  : in  std_logic                     := 'X';             -- readdatavalid
			dram_ctrl_s1_waitrequest                                    : in  std_logic                     := 'X';             -- waitrequest
			dram_ctrl_s1_chipselect                                     : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                           : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                            : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                      : out std_logic;                                        -- chipselect
			LCD_Controller_avalon_slave_0_address                       : out std_logic_vector(0 downto 0);                     -- address
			LCD_Controller_avalon_slave_0_write                         : out std_logic;                                        -- write
			LCD_Controller_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			LCD_Controller_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			LCD_Reset_N_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			LCD_Reset_N_s1_write                                        : out std_logic;                                        -- write
			LCD_Reset_N_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LCD_Reset_N_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			LCD_Reset_N_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Pitch_dummy_0_sp_address                                    : out std_logic_vector(1 downto 0);                     -- address
			Pitch_dummy_0_sp_write                                      : out std_logic;                                        -- write
			Pitch_dummy_0_sp_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pitch_dummy_0_sp_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			sysid_control_slave_address                                 : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_s1_address                                            : out std_logic_vector(2 downto 0);                     -- address
			timer_s1_write                                              : out std_logic;                                        -- write
			timer_s1_readdata                                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_s1_writedata                                          : out std_logic_vector(15 downto 0);                    -- writedata
			timer_s1_chipselect                                         : out std_logic;                                        -- chipselect
			touch_panel_busy_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			touch_panel_busy_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			touch_panel_pen_irq_n_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			touch_panel_pen_irq_n_s1_write                              : out std_logic;                                        -- write
			touch_panel_pen_irq_n_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			touch_panel_pen_irq_n_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			touch_panel_pen_irq_n_s1_chipselect                         : out std_logic;                                        -- chipselect
			touch_panel_spi_spi_control_port_address                    : out std_logic_vector(2 downto 0);                     -- address
			touch_panel_spi_spi_control_port_write                      : out std_logic;                                        -- write
			touch_panel_spi_spi_control_port_read                       : out std_logic;                                        -- read
			touch_panel_spi_spi_control_port_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			touch_panel_spi_spi_control_port_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			touch_panel_spi_spi_control_port_chipselect                 : out std_logic;                                        -- chipselect
			Volume_dummy_0_sp_address                                   : out std_logic_vector(0 downto 0);                     -- address
			Volume_dummy_0_sp_write                                     : out std_logic;                                        -- write
			Volume_dummy_0_sp_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Volume_dummy_0_sp_writedata                                 : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component system_mm_interconnect_0;

	component system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller;

	component system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component system_rst_controller_001;

	signal pll_outclk0_clk                                                               : std_logic;                     -- pll:outclk_0 -> [Pitch_dummy_0:csi_clk, Volume_dummy_0:csi_clk, cpu:clk, dram_ctrl:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, rst_controller_001:clk, sysid:clock, timer:clk]
	signal pll_outclk1_clk                                                               : std_logic;                     -- pll:outclk_1 -> [LCD_Controller:clk, LCD_Reset_N:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_0:pll_outclk1_clk, rst_controller:clk, touch_panel_busy:clk, touch_panel_pen_irq_n:clk, touch_panel_spi:clk]
	signal pll_outclk3_clk                                                               : std_logic;                     -- pll:outclk_3 -> [audio_and_video_config_0:clk, mm_interconnect_0:pll_outclk3_clk, rst_controller_002:clk]
	signal pll_outclk4_clk                                                               : std_logic;                     -- pll:outclk_4 -> [rst_controller_003:clk, ton_generation_dummy_0:clk]
	signal cpu_debug_reset_request_reset                                                 : std_logic;                     -- cpu:debug_reset_request -> [cpu_debug_reset_request_reset:in, mm_interconnect_0:dram_ctrl_reset_reset_bridge_in_reset_reset]
	signal cpu_data_master_readdata                                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                                   : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                       : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                    : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                          : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                                 : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                                         : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                     : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                                   : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                          : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect                    : std_logic;                     -- mm_interconnect_0:LCD_Controller_avalon_slave_0_chipselect -> mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:LCD_Controller_avalon_slave_0_address -> LCD_Controller:s_address
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_write                         : std_logic;                     -- mm_interconnect_0:LCD_Controller_avalon_slave_0_write -> mm_interconnect_0_lcd_controller_avalon_slave_0_write:in
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_Controller_avalon_slave_0_writedata -> LCD_Controller:s_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                                : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                                : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                             : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                             : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                    : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_dram_ctrl_s1_chipselect                                     : std_logic;                     -- mm_interconnect_0:dram_ctrl_s1_chipselect -> dram_ctrl:az_cs
	signal mm_interconnect_0_dram_ctrl_s1_readdata                                       : std_logic_vector(15 downto 0); -- dram_ctrl:za_data -> mm_interconnect_0:dram_ctrl_s1_readdata
	signal mm_interconnect_0_dram_ctrl_s1_waitrequest                                    : std_logic;                     -- dram_ctrl:za_waitrequest -> mm_interconnect_0:dram_ctrl_s1_waitrequest
	signal mm_interconnect_0_dram_ctrl_s1_address                                        : std_logic_vector(24 downto 0); -- mm_interconnect_0:dram_ctrl_s1_address -> dram_ctrl:az_addr
	signal mm_interconnect_0_dram_ctrl_s1_read                                           : std_logic;                     -- mm_interconnect_0:dram_ctrl_s1_read -> mm_interconnect_0_dram_ctrl_s1_read:in
	signal mm_interconnect_0_dram_ctrl_s1_byteenable                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:dram_ctrl_s1_byteenable -> mm_interconnect_0_dram_ctrl_s1_byteenable:in
	signal mm_interconnect_0_dram_ctrl_s1_readdatavalid                                  : std_logic;                     -- dram_ctrl:za_valid -> mm_interconnect_0:dram_ctrl_s1_readdatavalid
	signal mm_interconnect_0_dram_ctrl_s1_write                                          : std_logic;                     -- mm_interconnect_0:dram_ctrl_s1_write -> mm_interconnect_0_dram_ctrl_s1_write:in
	signal mm_interconnect_0_dram_ctrl_s1_writedata                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:dram_ctrl_s1_writedata -> dram_ctrl:az_data
	signal mm_interconnect_0_lcd_reset_n_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:LCD_Reset_N_s1_chipselect -> LCD_Reset_N:chipselect
	signal mm_interconnect_0_lcd_reset_n_s1_readdata                                     : std_logic_vector(31 downto 0); -- LCD_Reset_N:readdata -> mm_interconnect_0:LCD_Reset_N_s1_readdata
	signal mm_interconnect_0_lcd_reset_n_s1_address                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LCD_Reset_N_s1_address -> LCD_Reset_N:address
	signal mm_interconnect_0_lcd_reset_n_s1_write                                        : std_logic;                     -- mm_interconnect_0:LCD_Reset_N_s1_write -> mm_interconnect_0_lcd_reset_n_s1_write:in
	signal mm_interconnect_0_lcd_reset_n_s1_writedata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_Reset_N_s1_writedata -> LCD_Reset_N:writedata
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:touch_panel_pen_irq_n_s1_chipselect -> touch_panel_pen_irq_n:chipselect
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata                           : std_logic_vector(31 downto 0); -- touch_panel_pen_irq_n:readdata -> mm_interconnect_0:touch_panel_pen_irq_n_s1_readdata
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:touch_panel_pen_irq_n_s1_address -> touch_panel_pen_irq_n:address
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_write                              : std_logic;                     -- mm_interconnect_0:touch_panel_pen_irq_n_s1_write -> mm_interconnect_0_touch_panel_pen_irq_n_s1_write:in
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:touch_panel_pen_irq_n_s1_writedata -> touch_panel_pen_irq_n:writedata
	signal mm_interconnect_0_touch_panel_busy_s1_readdata                                : std_logic_vector(31 downto 0); -- touch_panel_busy:readdata -> mm_interconnect_0:touch_panel_busy_s1_readdata
	signal mm_interconnect_0_touch_panel_busy_s1_address                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:touch_panel_busy_s1_address -> touch_panel_busy:address
	signal mm_interconnect_0_timer_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	signal mm_interconnect_0_timer_s1_readdata                                           : std_logic_vector(15 downto 0); -- timer:readdata -> mm_interconnect_0:timer_s1_readdata
	signal mm_interconnect_0_timer_s1_address                                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_s1_address -> timer:address
	signal mm_interconnect_0_timer_s1_write                                              : std_logic;                     -- mm_interconnect_0:timer_s1_write -> mm_interconnect_0_timer_s1_write:in
	signal mm_interconnect_0_timer_s1_writedata                                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_s1_writedata -> timer:writedata
	signal mm_interconnect_0_pitch_dummy_0_sp_readdata                                   : std_logic_vector(31 downto 0); -- Pitch_dummy_0:avs_sP_readdata -> mm_interconnect_0:Pitch_dummy_0_sp_readdata
	signal mm_interconnect_0_pitch_dummy_0_sp_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Pitch_dummy_0_sp_address -> Pitch_dummy_0:avs_sP_address
	signal mm_interconnect_0_pitch_dummy_0_sp_write                                      : std_logic;                     -- mm_interconnect_0:Pitch_dummy_0_sp_write -> Pitch_dummy_0:avs_sP_write
	signal mm_interconnect_0_pitch_dummy_0_sp_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:Pitch_dummy_0_sp_writedata -> Pitch_dummy_0:avs_sP_writedata
	signal mm_interconnect_0_volume_dummy_0_sp_readdata                                  : std_logic_vector(31 downto 0); -- Volume_dummy_0:avs_sP_readdata -> mm_interconnect_0:Volume_dummy_0_sp_readdata
	signal mm_interconnect_0_volume_dummy_0_sp_address                                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:Volume_dummy_0_sp_address -> Volume_dummy_0:avs_sP_address
	signal mm_interconnect_0_volume_dummy_0_sp_write                                     : std_logic;                     -- mm_interconnect_0:Volume_dummy_0_sp_write -> Volume_dummy_0:avs_sP_write
	signal mm_interconnect_0_volume_dummy_0_sp_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:Volume_dummy_0_sp_writedata -> Volume_dummy_0:avs_sP_writedata
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect                 : std_logic;                     -- mm_interconnect_0:touch_panel_spi_spi_control_port_chipselect -> touch_panel_spi:spi_select
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_readdata                   : std_logic_vector(15 downto 0); -- touch_panel_spi:data_to_cpu -> mm_interconnect_0:touch_panel_spi_spi_control_port_readdata
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:touch_panel_spi_spi_control_port_address -> touch_panel_spi:mem_addr
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_read                       : std_logic;                     -- mm_interconnect_0:touch_panel_spi_spi_control_port_read -> mm_interconnect_0_touch_panel_spi_spi_control_port_read:in
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_write                      : std_logic;                     -- mm_interconnect_0:touch_panel_spi_spi_control_port_write -> mm_interconnect_0_touch_panel_spi_spi_control_port_write:in
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:touch_panel_spi_spi_control_port_writedata -> touch_panel_spi:data_from_cpu
	signal irq_mapper_receiver1_irq                                                      : std_logic;                     -- timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver3_irq                                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal irq_mapper_receiver0_irq                                                      : std_logic;                     -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                                 : std_logic_vector(0 downto 0);  -- touch_panel_pen_irq_n:irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver2_irq                                                      : std_logic;                     -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_001_receiver_irq                                             : std_logic_vector(0 downto 0);  -- touch_panel_spi:irq -> irq_synchronizer_001:receiver_irq
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_interconnect_0:LCD_Controller_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                            : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                                        : std_logic;                     -- rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                                            : std_logic;                     -- rst_controller_002:reset_out -> [audio_and_video_config_0:reset, mm_interconnect_0:audio_and_video_config_0_reset_reset_bridge_in_reset_reset]
	signal rst_controller_003_reset_out_reset                                            : std_logic;                     -- rst_controller_003:reset_out -> rst_controller_003_reset_out_reset:in
	signal reset_reset_n_ports_inv                                                       : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal cpu_debug_reset_request_reset_ports_inv                                       : std_logic;                     -- cpu_debug_reset_request_reset:inv -> dram_ctrl:reset_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv                  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect_ports_inv          : std_logic;                     -- mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect:inv -> LCD_Controller:s_chipselect_n
	signal mm_interconnect_0_lcd_controller_avalon_slave_0_write_ports_inv               : std_logic;                     -- mm_interconnect_0_lcd_controller_avalon_slave_0_write:inv -> LCD_Controller:s_write_n
	signal mm_interconnect_0_dram_ctrl_s1_read_ports_inv                                 : std_logic;                     -- mm_interconnect_0_dram_ctrl_s1_read:inv -> dram_ctrl:az_rd_n
	signal mm_interconnect_0_dram_ctrl_s1_byteenable_ports_inv                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0_dram_ctrl_s1_byteenable:inv -> dram_ctrl:az_be_n
	signal mm_interconnect_0_dram_ctrl_s1_write_ports_inv                                : std_logic;                     -- mm_interconnect_0_dram_ctrl_s1_write:inv -> dram_ctrl:az_wr_n
	signal mm_interconnect_0_lcd_reset_n_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_lcd_reset_n_s1_write:inv -> LCD_Reset_N:write_n
	signal mm_interconnect_0_touch_panel_pen_irq_n_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_touch_panel_pen_irq_n_s1_write:inv -> touch_panel_pen_irq_n:write_n
	signal mm_interconnect_0_timer_s1_write_ports_inv                                    : std_logic;                     -- mm_interconnect_0_timer_s1_write:inv -> timer:write_n
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_read_ports_inv             : std_logic;                     -- mm_interconnect_0_touch_panel_spi_spi_control_port_read:inv -> touch_panel_spi:read_n
	signal mm_interconnect_0_touch_panel_spi_spi_control_port_write_ports_inv            : std_logic;                     -- mm_interconnect_0_touch_panel_spi_spi_control_port_write:inv -> touch_panel_spi:write_n
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [LCD_Controller:reset_n, LCD_Reset_N:reset_n, touch_panel_busy:reset_n, touch_panel_pen_irq_n:reset_n, touch_panel_spi:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [Pitch_dummy_0:rsi_reset_n, Volume_dummy_0:rsi_reset_n, cpu:reset_n, jtag_uart:rst_n, sysid:reset_n, timer:reset_n]
	signal rst_controller_003_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> ton_generation_dummy_0:reset_n

begin

	lcd_controller : component LT24_Controller
		port map (
			clk            => pll_outclk1_clk,                                                      --          clock.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                             --          reset.reset_n
			s_chipselect_n => mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			s_write_n      => mm_interconnect_0_lcd_controller_avalon_slave_0_write_ports_inv,      --               .write_n
			s_writedata    => mm_interconnect_0_lcd_controller_avalon_slave_0_writedata,            --               .writedata
			s_address      => mm_interconnect_0_lcd_controller_avalon_slave_0_address(0),           --               .address
			lt24_cs        => lcd_controller_conduit_end_lt24_cs,                                   --    conduit_end.lt24_cs
			lt24_data      => lcd_controller_conduit_end_lt24_data,                                 --               .lt24_data
			lt24_rd        => lcd_controller_conduit_end_lt24_rd,                                   --               .lt24_rd
			lt24_wr        => lcd_controller_conduit_end_lt24_wr,                                   --               .lt24_wr
			lt24_rs        => lcd_controller_conduit_end_lt24_rs                                    --               .lt24_rs
		);

	lcd_reset_n : component system_LCD_Reset_N
		port map (
			clk        => pll_outclk1_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_lcd_reset_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_lcd_reset_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_lcd_reset_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_lcd_reset_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_lcd_reset_n_s1_readdata,        --                    .readdata
			out_port   => lcd_reset_n_external_connection_export            -- external_connection.export
		);

	pitch_dummy_0 : component pitch_dummy
		generic map (
			dat_len_avl => 31,
			data_freq   => "00000000000000001111101000000000",
			data_freq1  => "00000000000000000111110100000000"
		)
		port map (
			avs_sP_address   => mm_interconnect_0_pitch_dummy_0_sp_address,   --            sp.address
			avs_sP_readdata  => mm_interconnect_0_pitch_dummy_0_sp_readdata,  --              .readdata
			avs_sP_write     => mm_interconnect_0_pitch_dummy_0_sp_write,     --              .write
			avs_sP_writedata => mm_interconnect_0_pitch_dummy_0_sp_writedata, --              .writedata
			coe_led_gli      => led_gli_export,                               -- conduit_end_0.export
			rsi_reset_n      => rst_controller_001_reset_out_reset_ports_inv, --         reset.reset_n
			csi_clk          => pll_outclk0_clk,                              --         clock.clk
			coe_led_delay    => led_delay_export                              --   conduit_end.export
		);

	volume_dummy_0 : component volume_dummy
		generic map (
			dat_len_avl => 31,
			data_freq   => "00000000000000001111101000000000",
			data_freq1  => "00000000000000000111110100000000"
		)
		port map (
			avs_sP_address   => mm_interconnect_0_volume_dummy_0_sp_address(0), --            sp.address
			avs_sP_readdata  => mm_interconnect_0_volume_dummy_0_sp_readdata,   --              .readdata
			avs_sP_write     => mm_interconnect_0_volume_dummy_0_sp_write,      --              .write
			avs_sP_writedata => mm_interconnect_0_volume_dummy_0_sp_writedata,  --              .writedata
			coe_led_vol      => led_vol_export,                                 -- conduit_end_0.export
			rsi_reset_n      => rst_controller_001_reset_out_reset_ports_inv,   --         reset.reset_n
			csi_clk          => pll_outclk0_clk                                 --         clock.clk
		);

	audio_and_video_config_0 : component system_audio_and_video_config_0
		port map (
			clk         => pll_outclk3_clk,                                                               --                    clk.clk
			reset       => rst_controller_002_reset_out_reset,                                            --                  reset.reset
			address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_and_video_config_0_external_interface_SDAT,                              --     external_interface.export
			I2C_SCLK    => audio_and_video_config_0_external_interface_SCLK                               --                       .export
		);

	cpu : component system_cpu
		port map (
			clk                                 => pll_outclk0_clk,                                   --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	dram_ctrl : component system_dram_ctrl
		port map (
			clk            => pll_outclk0_clk,                                     --   clk.clk
			reset_n        => cpu_debug_reset_request_reset_ports_inv,             -- reset.reset_n
			az_addr        => mm_interconnect_0_dram_ctrl_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_dram_ctrl_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_dram_ctrl_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_dram_ctrl_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_dram_ctrl_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_dram_ctrl_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_dram_ctrl_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_dram_ctrl_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_dram_ctrl_s1_waitrequest,          --      .waitrequest
			zs_addr        => dram_ctrl_wire_addr,                                 --  wire.export
			zs_ba          => dram_ctrl_wire_ba,                                   --      .export
			zs_cas_n       => dram_ctrl_wire_cas_n,                                --      .export
			zs_cke         => dram_ctrl_wire_cke,                                  --      .export
			zs_cs_n        => dram_ctrl_wire_cs_n,                                 --      .export
			zs_dq          => dram_ctrl_wire_dq,                                   --      .export
			zs_dqm         => dram_ctrl_wire_dqm,                                  --      .export
			zs_ras_n       => dram_ctrl_wire_ras_n,                                --      .export
			zs_we_n        => dram_ctrl_wire_we_n                                  --      .export
		);

	jtag_uart : component system_jtag_uart
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver3_irq                                       --               irq.irq
		);

	pll : component system_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => pll_outclk1_clk,         -- outclk1.clk
			outclk_2 => sdram_clk_clk,           -- outclk2.clk
			outclk_3 => pll_outclk3_clk,         -- outclk3.clk
			outclk_4 => pll_outclk4_clk,         -- outclk4.clk
			outclk_5 => aud_xck_clk,             -- outclk5.clk
			locked   => open                     -- (terminated)
		);

	sysid : component system_sysid
		port map (
			clock    => pll_outclk0_clk,                                  --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer : component system_timer
		port map (
			clk        => pll_outclk0_clk,                              --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_s1_address,           --    s1.address
			writedata  => mm_interconnect_0_timer_s1_writedata,         --      .writedata
			readdata   => mm_interconnect_0_timer_s1_readdata,          --      .readdata
			chipselect => mm_interconnect_0_timer_s1_chipselect,        --      .chipselect
			write_n    => mm_interconnect_0_timer_s1_write_ports_inv,   --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	ton_generation_dummy_0 : component sine1kHz
		port map (
			reset_n          => rst_controller_003_reset_out_reset_ports_inv, --         reset.reset_n
			clk              => pll_outclk4_clk,                              --         clock.clk
			coe_AUD2_DACDAT  => dacdat_export,                                -- conduit_end_0.export
			coe_AUD1_BCLK    => bclk_export,                                  --   conduit_end.export
			coe_AUD3_DACLRCK => daclrck_export                                -- conduit_end_1.export
		);

	touch_panel_busy : component system_touch_panel_busy
		port map (
			clk      => pll_outclk1_clk,                                --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address  => mm_interconnect_0_touch_panel_busy_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_touch_panel_busy_s1_readdata, --                    .readdata
			in_port  => touch_panel_busy_external_connection_export     -- external_connection.export
		);

	touch_panel_pen_irq_n : component system_touch_panel_pen_irq_n
		port map (
			clk        => pll_outclk1_clk,                                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => mm_interconnect_0_touch_panel_pen_irq_n_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_touch_panel_pen_irq_n_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata,        --                    .readdata
			in_port    => touch_panel_pen_irq_n_external_connection_export,           -- external_connection.export
			irq        => irq_synchronizer_receiver_irq(0)                            --                 irq.irq
		);

	touch_panel_spi : component system_touch_panel_spi
		port map (
			clk           => pll_outclk1_clk,                                                    --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                           --            reset.reset_n
			data_from_cpu => mm_interconnect_0_touch_panel_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_touch_panel_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_touch_panel_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_touch_panel_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_touch_panel_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_synchronizer_001_receiver_irq(0),                               --              irq.irq
			MISO          => touch_panel_spi_external_MISO,                                      --         external.export
			MOSI          => touch_panel_spi_external_MOSI,                                      --                 .export
			SCLK          => touch_panel_spi_external_SCLK,                                      --                 .export
			SS_n          => touch_panel_spi_external_SS_n                                       --                 .export
		);

	mm_interconnect_0 : component system_mm_interconnect_0
		port map (
			pll_outclk0_clk                                             => pll_outclk0_clk,                                                               --                                          pll_outclk0.clk
			pll_outclk1_clk                                             => pll_outclk1_clk,                                                               --                                          pll_outclk1.clk
			pll_outclk3_clk                                             => pll_outclk3_clk,                                                               --                                          pll_outclk3.clk
			audio_and_video_config_0_reset_reset_bridge_in_reset_reset  => rst_controller_002_reset_out_reset,                                            -- audio_and_video_config_0_reset_reset_bridge_in_reset.reset
			cpu_reset_reset_bridge_in_reset_reset                       => rst_controller_001_reset_out_reset,                                            --                      cpu_reset_reset_bridge_in_reset.reset
			dram_ctrl_reset_reset_bridge_in_reset_reset                 => cpu_debug_reset_request_reset,                                                 --                dram_ctrl_reset_reset_bridge_in_reset.reset
			LCD_Controller_reset_reset_bridge_in_reset_reset            => rst_controller_reset_out_reset,                                                --           LCD_Controller_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                     => cpu_data_master_address,                                                       --                                      cpu_data_master.address
			cpu_data_master_waitrequest                                 => cpu_data_master_waitrequest,                                                   --                                                     .waitrequest
			cpu_data_master_byteenable                                  => cpu_data_master_byteenable,                                                    --                                                     .byteenable
			cpu_data_master_read                                        => cpu_data_master_read,                                                          --                                                     .read
			cpu_data_master_readdata                                    => cpu_data_master_readdata,                                                      --                                                     .readdata
			cpu_data_master_readdatavalid                               => cpu_data_master_readdatavalid,                                                 --                                                     .readdatavalid
			cpu_data_master_write                                       => cpu_data_master_write,                                                         --                                                     .write
			cpu_data_master_writedata                                   => cpu_data_master_writedata,                                                     --                                                     .writedata
			cpu_data_master_debugaccess                                 => cpu_data_master_debugaccess,                                                   --                                                     .debugaccess
			cpu_instruction_master_address                              => cpu_instruction_master_address,                                                --                               cpu_instruction_master.address
			cpu_instruction_master_waitrequest                          => cpu_instruction_master_waitrequest,                                            --                                                     .waitrequest
			cpu_instruction_master_read                                 => cpu_instruction_master_read,                                                   --                                                     .read
			cpu_instruction_master_readdata                             => cpu_instruction_master_readdata,                                               --                                                     .readdata
			cpu_instruction_master_readdatavalid                        => cpu_instruction_master_readdatavalid,                                          --                                                     .readdatavalid
			audio_and_video_config_0_avalon_av_config_slave_address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     --      audio_and_video_config_0_avalon_av_config_slave.address
			audio_and_video_config_0_avalon_av_config_slave_write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                                                     .write
			audio_and_video_config_0_avalon_av_config_slave_read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                                                     .read
			audio_and_video_config_0_avalon_av_config_slave_readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                                                     .readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                                                     .writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                                                     .byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                                                     .waitrequest
			cpu_debug_mem_slave_address                                 => mm_interconnect_0_cpu_debug_mem_slave_address,                                 --                                  cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                   => mm_interconnect_0_cpu_debug_mem_slave_write,                                   --                                                     .write
			cpu_debug_mem_slave_read                                    => mm_interconnect_0_cpu_debug_mem_slave_read,                                    --                                                     .read
			cpu_debug_mem_slave_readdata                                => mm_interconnect_0_cpu_debug_mem_slave_readdata,                                --                                                     .readdata
			cpu_debug_mem_slave_writedata                               => mm_interconnect_0_cpu_debug_mem_slave_writedata,                               --                                                     .writedata
			cpu_debug_mem_slave_byteenable                              => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                              --                                                     .byteenable
			cpu_debug_mem_slave_waitrequest                             => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                             --                                                     .waitrequest
			cpu_debug_mem_slave_debugaccess                             => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                             --                                                     .debugaccess
			dram_ctrl_s1_address                                        => mm_interconnect_0_dram_ctrl_s1_address,                                        --                                         dram_ctrl_s1.address
			dram_ctrl_s1_write                                          => mm_interconnect_0_dram_ctrl_s1_write,                                          --                                                     .write
			dram_ctrl_s1_read                                           => mm_interconnect_0_dram_ctrl_s1_read,                                           --                                                     .read
			dram_ctrl_s1_readdata                                       => mm_interconnect_0_dram_ctrl_s1_readdata,                                       --                                                     .readdata
			dram_ctrl_s1_writedata                                      => mm_interconnect_0_dram_ctrl_s1_writedata,                                      --                                                     .writedata
			dram_ctrl_s1_byteenable                                     => mm_interconnect_0_dram_ctrl_s1_byteenable,                                     --                                                     .byteenable
			dram_ctrl_s1_readdatavalid                                  => mm_interconnect_0_dram_ctrl_s1_readdatavalid,                                  --                                                     .readdatavalid
			dram_ctrl_s1_waitrequest                                    => mm_interconnect_0_dram_ctrl_s1_waitrequest,                                    --                                                     .waitrequest
			dram_ctrl_s1_chipselect                                     => mm_interconnect_0_dram_ctrl_s1_chipselect,                                     --                                                     .chipselect
			jtag_uart_avalon_jtag_slave_address                         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,                         --                          jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,                           --                                                     .write
			jtag_uart_avalon_jtag_slave_read                            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                            --                                                     .read
			jtag_uart_avalon_jtag_slave_readdata                        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,                        --                                                     .readdata
			jtag_uart_avalon_jtag_slave_writedata                       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,                       --                                                     .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,                     --                                                     .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,                      --                                                     .chipselect
			LCD_Controller_avalon_slave_0_address                       => mm_interconnect_0_lcd_controller_avalon_slave_0_address,                       --                        LCD_Controller_avalon_slave_0.address
			LCD_Controller_avalon_slave_0_write                         => mm_interconnect_0_lcd_controller_avalon_slave_0_write,                         --                                                     .write
			LCD_Controller_avalon_slave_0_writedata                     => mm_interconnect_0_lcd_controller_avalon_slave_0_writedata,                     --                                                     .writedata
			LCD_Controller_avalon_slave_0_chipselect                    => mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect,                    --                                                     .chipselect
			LCD_Reset_N_s1_address                                      => mm_interconnect_0_lcd_reset_n_s1_address,                                      --                                       LCD_Reset_N_s1.address
			LCD_Reset_N_s1_write                                        => mm_interconnect_0_lcd_reset_n_s1_write,                                        --                                                     .write
			LCD_Reset_N_s1_readdata                                     => mm_interconnect_0_lcd_reset_n_s1_readdata,                                     --                                                     .readdata
			LCD_Reset_N_s1_writedata                                    => mm_interconnect_0_lcd_reset_n_s1_writedata,                                    --                                                     .writedata
			LCD_Reset_N_s1_chipselect                                   => mm_interconnect_0_lcd_reset_n_s1_chipselect,                                   --                                                     .chipselect
			Pitch_dummy_0_sp_address                                    => mm_interconnect_0_pitch_dummy_0_sp_address,                                    --                                     Pitch_dummy_0_sp.address
			Pitch_dummy_0_sp_write                                      => mm_interconnect_0_pitch_dummy_0_sp_write,                                      --                                                     .write
			Pitch_dummy_0_sp_readdata                                   => mm_interconnect_0_pitch_dummy_0_sp_readdata,                                   --                                                     .readdata
			Pitch_dummy_0_sp_writedata                                  => mm_interconnect_0_pitch_dummy_0_sp_writedata,                                  --                                                     .writedata
			sysid_control_slave_address                                 => mm_interconnect_0_sysid_control_slave_address,                                 --                                  sysid_control_slave.address
			sysid_control_slave_readdata                                => mm_interconnect_0_sysid_control_slave_readdata,                                --                                                     .readdata
			timer_s1_address                                            => mm_interconnect_0_timer_s1_address,                                            --                                             timer_s1.address
			timer_s1_write                                              => mm_interconnect_0_timer_s1_write,                                              --                                                     .write
			timer_s1_readdata                                           => mm_interconnect_0_timer_s1_readdata,                                           --                                                     .readdata
			timer_s1_writedata                                          => mm_interconnect_0_timer_s1_writedata,                                          --                                                     .writedata
			timer_s1_chipselect                                         => mm_interconnect_0_timer_s1_chipselect,                                         --                                                     .chipselect
			touch_panel_busy_s1_address                                 => mm_interconnect_0_touch_panel_busy_s1_address,                                 --                                  touch_panel_busy_s1.address
			touch_panel_busy_s1_readdata                                => mm_interconnect_0_touch_panel_busy_s1_readdata,                                --                                                     .readdata
			touch_panel_pen_irq_n_s1_address                            => mm_interconnect_0_touch_panel_pen_irq_n_s1_address,                            --                             touch_panel_pen_irq_n_s1.address
			touch_panel_pen_irq_n_s1_write                              => mm_interconnect_0_touch_panel_pen_irq_n_s1_write,                              --                                                     .write
			touch_panel_pen_irq_n_s1_readdata                           => mm_interconnect_0_touch_panel_pen_irq_n_s1_readdata,                           --                                                     .readdata
			touch_panel_pen_irq_n_s1_writedata                          => mm_interconnect_0_touch_panel_pen_irq_n_s1_writedata,                          --                                                     .writedata
			touch_panel_pen_irq_n_s1_chipselect                         => mm_interconnect_0_touch_panel_pen_irq_n_s1_chipselect,                         --                                                     .chipselect
			touch_panel_spi_spi_control_port_address                    => mm_interconnect_0_touch_panel_spi_spi_control_port_address,                    --                     touch_panel_spi_spi_control_port.address
			touch_panel_spi_spi_control_port_write                      => mm_interconnect_0_touch_panel_spi_spi_control_port_write,                      --                                                     .write
			touch_panel_spi_spi_control_port_read                       => mm_interconnect_0_touch_panel_spi_spi_control_port_read,                       --                                                     .read
			touch_panel_spi_spi_control_port_readdata                   => mm_interconnect_0_touch_panel_spi_spi_control_port_readdata,                   --                                                     .readdata
			touch_panel_spi_spi_control_port_writedata                  => mm_interconnect_0_touch_panel_spi_spi_control_port_writedata,                  --                                                     .writedata
			touch_panel_spi_spi_control_port_chipselect                 => mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect,                 --                                                     .chipselect
			Volume_dummy_0_sp_address                                   => mm_interconnect_0_volume_dummy_0_sp_address,                                   --                                    Volume_dummy_0_sp.address
			Volume_dummy_0_sp_write                                     => mm_interconnect_0_volume_dummy_0_sp_write,                                     --                                                     .write
			Volume_dummy_0_sp_readdata                                  => mm_interconnect_0_volume_dummy_0_sp_readdata,                                  --                                                     .readdata
			Volume_dummy_0_sp_writedata                                 => mm_interconnect_0_volume_dummy_0_sp_writedata                                  --                                                     .writedata
		);

	irq_mapper : component system_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                    --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk1_clk,                    --       receiver_clk.clk
			sender_clk     => pll_outclk0_clk,                    --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => pll_outclk1_clk,                    --       receiver_clk.clk
			sender_clk     => pll_outclk0_clk,                    --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	rst_controller : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => pll_outclk1_clk,                --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_outclk0_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_outclk3_clk,                    --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_outclk4_clk,                    --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	cpu_debug_reset_request_reset_ports_inv <= not cpu_debug_reset_request_reset;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_lcd_controller_avalon_slave_0_chipselect;

	mm_interconnect_0_lcd_controller_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_lcd_controller_avalon_slave_0_write;

	mm_interconnect_0_dram_ctrl_s1_read_ports_inv <= not mm_interconnect_0_dram_ctrl_s1_read;

	mm_interconnect_0_dram_ctrl_s1_byteenable_ports_inv <= not mm_interconnect_0_dram_ctrl_s1_byteenable;

	mm_interconnect_0_dram_ctrl_s1_write_ports_inv <= not mm_interconnect_0_dram_ctrl_s1_write;

	mm_interconnect_0_lcd_reset_n_s1_write_ports_inv <= not mm_interconnect_0_lcd_reset_n_s1_write;

	mm_interconnect_0_touch_panel_pen_irq_n_s1_write_ports_inv <= not mm_interconnect_0_touch_panel_pen_irq_n_s1_write;

	mm_interconnect_0_timer_s1_write_ports_inv <= not mm_interconnect_0_timer_s1_write;

	mm_interconnect_0_touch_panel_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_touch_panel_spi_spi_control_port_read;

	mm_interconnect_0_touch_panel_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_touch_panel_spi_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of system
