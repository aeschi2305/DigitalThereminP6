-- altera_asmi_parallel_digital_theremin_epcq_controller_0.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity altera_asmi_parallel_digital_theremin_epcq_controller_0 is
	port (
		clkin          : in  std_logic                     := '0';             --          clkin.clk
		fast_read      : in  std_logic                     := '0';             --      fast_read.fast_read
		rden           : in  std_logic                     := '0';             --           rden.rden
		addr           : in  std_logic_vector(23 downto 0) := (others => '0'); --           addr.addr
		read_status    : in  std_logic                     := '0';             --    read_status.read_status
		write          : in  std_logic                     := '0';             --          write.write
		datain         : in  std_logic_vector(7 downto 0)  := (others => '0'); --         datain.datain
		shift_bytes    : in  std_logic                     := '0';             --    shift_bytes.shift_bytes
		sector_protect : in  std_logic                     := '0';             -- sector_protect.sector_protect
		sector_erase   : in  std_logic                     := '0';             --   sector_erase.sector_erase
		bulk_erase     : in  std_logic                     := '0';             --     bulk_erase.bulk_erase
		wren           : in  std_logic                     := '0';             --           wren.wren
		read_rdid      : in  std_logic                     := '0';             --      read_rdid.read_rdid
		reset          : in  std_logic                     := '0';             --          reset.reset
		read_dummyclk  : in  std_logic                     := '0';             --  read_dummyclk.read_dummyclk
		dataout        : out std_logic_vector(7 downto 0);                     --        dataout.dataout
		busy           : out std_logic;                                        --           busy.busy
		data_valid     : out std_logic;                                        --     data_valid.data_valid
		status_out     : out std_logic_vector(7 downto 0);                     --     status_out.status_out
		illegal_write  : out std_logic;                                        --  illegal_write.illegal_write
		illegal_erase  : out std_logic;                                        --  illegal_erase.illegal_erase
		rdid_out       : out std_logic_vector(7 downto 0)                      --       rdid_out.rdid_out
	);
end entity altera_asmi_parallel_digital_theremin_epcq_controller_0;

architecture rtl of altera_asmi_parallel_digital_theremin_epcq_controller_0 is
	component digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0 is
		port (
			clkin          : in  std_logic                     := 'X';             -- clk
			fast_read      : in  std_logic                     := 'X';             -- fast_read
			rden           : in  std_logic                     := 'X';             -- rden
			addr           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- addr
			read_status    : in  std_logic                     := 'X';             -- read_status
			write          : in  std_logic                     := 'X';             -- write
			datain         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- datain
			shift_bytes    : in  std_logic                     := 'X';             -- shift_bytes
			sector_protect : in  std_logic                     := 'X';             -- sector_protect
			sector_erase   : in  std_logic                     := 'X';             -- sector_erase
			bulk_erase     : in  std_logic                     := 'X';             -- bulk_erase
			wren           : in  std_logic                     := 'X';             -- wren
			read_rdid      : in  std_logic                     := 'X';             -- read_rdid
			reset          : in  std_logic                     := 'X';             -- reset
			read_dummyclk  : in  std_logic                     := 'X';             -- read_dummyclk
			dataout        : out std_logic_vector(7 downto 0);                     -- dataout
			busy           : out std_logic;                                        -- busy
			data_valid     : out std_logic;                                        -- data_valid
			status_out     : out std_logic_vector(7 downto 0);                     -- status_out
			illegal_write  : out std_logic;                                        -- illegal_write
			illegal_erase  : out std_logic;                                        -- illegal_erase
			rdid_out       : out std_logic_vector(7 downto 0)                      -- rdid_out
		);
	end component digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0;

begin

	altera_asmi_parallel_digital_theremin_epcq_controller_0 : component digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0_altera_asmi_parallel_digital_theremin_epcq_controller_0
		port map (
			clkin          => clkin,          --          clkin.clk
			fast_read      => fast_read,      --      fast_read.fast_read
			rden           => rden,           --           rden.rden
			addr           => addr,           --           addr.addr
			read_status    => read_status,    --    read_status.read_status
			write          => write,          --          write.write
			datain         => datain,         --         datain.datain
			shift_bytes    => shift_bytes,    --    shift_bytes.shift_bytes
			sector_protect => sector_protect, -- sector_protect.sector_protect
			sector_erase   => sector_erase,   --   sector_erase.sector_erase
			bulk_erase     => bulk_erase,     --     bulk_erase.bulk_erase
			wren           => wren,           --           wren.wren
			read_rdid      => read_rdid,      --      read_rdid.read_rdid
			reset          => reset,          --          reset.reset
			read_dummyclk  => read_dummyclk,  --  read_dummyclk.read_dummyclk
			dataout        => dataout,        --        dataout.dataout
			busy           => busy,           --           busy.busy
			data_valid     => data_valid,     --     data_valid.data_valid
			status_out     => status_out,     --     status_out.status_out
			illegal_write  => illegal_write,  --  illegal_write.illegal_write
			illegal_erase  => illegal_erase,  --  illegal_erase.illegal_erase
			rdid_out       => rdid_out        --       rdid_out.rdid_out
		);

end architecture rtl; -- of altera_asmi_parallel_digital_theremin_epcq_controller_0
